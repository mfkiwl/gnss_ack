module gps_ack
(
	input wire clk,
	input wire rst,
	input wire i_sample,
	input wire [5:0] satelite,
	input wire [9:0] chip_delay,
	input wire [31:0] doppler,
	output wire [15:0] integrator
);








endmodule
